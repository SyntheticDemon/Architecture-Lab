library verilog;
use verilog.vl_types.all;
entity instruction_memory_tb is
end instruction_memory_tb;
