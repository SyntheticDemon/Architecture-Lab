library verilog;
use verilog.vl_types.all;
entity IF_Stage_Testbench is
end IF_Stage_Testbench;
