module moduleName (
    ports
);
    
endmodule